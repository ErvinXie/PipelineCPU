module WriteMem();






endmodule