module FetchInst(
    input clk,
    input rst
);



endmodule