module InstDecode();


endmodule