module WriteBack();


endmodule