`timescale 1ns / 1ps
`include "Marco.v"

module Imem(input clk,
            input rst,
            input[31:0] iaddr,
            output [31:0] idata);
    
    reg[31:0] mem[`IMEM_SIZE/4-1:0];
    
    wire[`IMEM_ADDR_WIDTH-1:0] addr;
    assign addr  = iaddr[`IMEM_ADDR_WIDTH-1:0];
    assign idata = mem[(addr>>2)];
    integer i;

    always@(negedge rst)begin

        mem[0]<=32'h3c180007;
        mem[1]<=32'h3c190008;
        mem[2]<=32'h24100140;
        mem[3]<=32'h241100f0;
        mem[4]<=32'h2412000e;
        mem[5]<=32'h2413000e;
        mem[6]<=32'h00121021;
        mem[7]<=32'h00131821;
        mem[8]<=32'h00122021;
        mem[9]<=32'h00022021;
        mem[10]<=32'h00032821;
        mem[11]<=32'h00023021;
        mem[12]<=32'h00063022;
        mem[13]<=32'h0c100019;
        mem[14]<=32'h00000000;
        mem[15]<=32'haf070000;
        mem[16]<=32'haf270000;
        mem[17]<=32'h26730001;
        mem[18]<=32'h1671fff3;
        mem[19]<=32'h00000000;
        mem[20]<=32'h26520001;
        mem[21]<=32'h1650ffef;
        mem[22]<=32'h00000000;
        mem[23]<=32'h08100028;
        mem[24]<=32'h00000000;
        mem[25]<=32'h3084000f;
        mem[26]<=32'h00042200;
        mem[27]<=32'h30a5000f;
        mem[28]<=32'h00052900;
        mem[29]<=32'h30c6000f;
        mem[30]<=32'h304203ff;
        mem[31]<=32'h00021300;
        mem[32]<=32'h306303ff;
        mem[33]<=32'h00031d80;
        mem[34]<=32'h00431025;
        mem[35]<=32'h00852025;
        mem[36]<=32'h00823825;
        mem[37]<=32'h00e63825;
        mem[38]<=32'h03e00008;
        mem[39]<=32'h00000000;
        mem[40]<=32'h00000000;
        mem[41]<=32'h00000000;
        mem[42]<=32'h00000000;
        mem[43]<=32'h00000000;
        mem[44]<=32'h00000000;
        mem[45]<=32'h00000000;
        mem[46]<=32'h00000000;
        mem[47]<=32'h00000000;
        mem[48]<=32'h00000000;
        mem[49]<=32'h00000000;
        mem[50]<=32'h00000000;
        mem[51]<=32'h00000000;
        mem[52]<=32'h00000000;
        mem[53]<=32'h00000000;
        mem[54]<=32'h00000000;
        mem[55]<=32'h00000000;
        mem[56]<=32'h00000000;
        mem[57]<=32'h00000000;
        mem[58]<=32'h00000000;
        mem[59]<=32'h00000000;
        mem[60]<=32'h00000000;
        mem[61]<=32'h00000000;
        mem[62]<=32'h00000000;
        mem[63]<=32'h00000000;
        mem[64]<=32'h00000000;
        mem[65]<=32'h00000000;
        mem[66]<=32'h00000000;
        mem[67]<=32'h00000000;
        mem[68]<=32'h00000000;
        mem[69]<=32'h00000000;
        mem[70]<=32'h00000000;
        mem[71]<=32'h00000000;
        mem[72]<=32'h00000000;
        mem[73]<=32'h00000000;
        mem[74]<=32'h00000000;
        mem[75]<=32'h00000000;
        mem[76]<=32'h00000000;
        mem[77]<=32'h00000000;
        mem[78]<=32'h00000000;
        mem[79]<=32'h00000000;
        mem[80]<=32'h00000000;
        mem[81]<=32'h00000000;
        mem[82]<=32'h00000000;
        mem[83]<=32'h00000000;
        mem[84]<=32'h00000000;
        mem[85]<=32'h00000000;
        mem[86]<=32'h00000000;
        mem[87]<=32'h00000000;
        mem[88]<=32'h00000000;
        mem[89]<=32'h00000000;
        mem[90]<=32'h00000000;
        mem[91]<=32'h00000000;
        mem[92]<=32'h00000000;
        mem[93]<=32'h00000000;
        mem[94]<=32'h00000000;
        mem[95]<=32'h00000000;
        mem[96]<=32'h00000000;
        mem[97]<=32'h00000000;
        mem[98]<=32'h00000000;
        mem[99]<=32'h00000000;
        mem[100]<=32'h00000000;
        mem[101]<=32'h00000000;
        mem[102]<=32'h00000000;
        mem[103]<=32'h00000000;
        mem[104]<=32'h00000000;
        mem[105]<=32'h00000000;
        mem[106]<=32'h00000000;
        mem[107]<=32'h00000000;
        mem[108]<=32'h00000000;
        mem[109]<=32'h00000000;
        mem[110]<=32'h00000000;
        mem[111]<=32'h00000000;
        mem[112]<=32'h00000000;
        mem[113]<=32'h00000000;
        mem[114]<=32'h00000000;
        mem[115]<=32'h00000000;
        mem[116]<=32'h00000000;
        mem[117]<=32'h00000000;
        mem[118]<=32'h00000000;
        mem[119]<=32'h00000000;
        mem[120]<=32'h00000000;
        mem[121]<=32'h00000000;
        mem[122]<=32'h00000000;
        mem[123]<=32'h00000000;
        mem[124]<=32'h00000000;
        mem[125]<=32'h00000000;
        mem[126]<=32'h00000000;
        mem[127]<=32'h00000000;
        mem[128]<=32'h00000000;
        mem[129]<=32'h00000000;
        mem[130]<=32'h00000000;
        mem[131]<=32'h00000000;
        mem[132]<=32'h00000000;
        mem[133]<=32'h00000000;
        mem[134]<=32'h00000000;
        mem[135]<=32'h00000000;
        mem[136]<=32'h00000000;
        mem[137]<=32'h00000000;
        mem[138]<=32'h00000000;
        mem[139]<=32'h00000000;
        mem[140]<=32'h00000000;
        mem[141]<=32'h00000000;
        mem[142]<=32'h00000000;
        mem[143]<=32'h00000000;
        mem[144]<=32'h00000000;
        mem[145]<=32'h00000000;
        mem[146]<=32'h00000000;
        mem[147]<=32'h00000000;
        mem[148]<=32'h00000000;
        mem[149]<=32'h00000000;
        mem[150]<=32'h00000000;
        mem[151]<=32'h00000000;
        mem[152]<=32'h00000000;
        mem[153]<=32'h00000000;
        mem[154]<=32'h00000000;
        mem[155]<=32'h00000000;
        mem[156]<=32'h00000000;
        mem[157]<=32'h00000000;
        mem[158]<=32'h00000000;
        mem[159]<=32'h00000000;
        mem[160]<=32'h00000000;
        mem[161]<=32'h00000000;
        mem[162]<=32'h00000000;
        mem[163]<=32'h00000000;
        mem[164]<=32'h00000000;
        mem[165]<=32'h00000000;
        mem[166]<=32'h00000000;
        mem[167]<=32'h00000000;
        mem[168]<=32'h00000000;
        mem[169]<=32'h00000000;
        mem[170]<=32'h00000000;
        mem[171]<=32'h00000000;
        mem[172]<=32'h00000000;
        mem[173]<=32'h00000000;
        mem[174]<=32'h00000000;
        mem[175]<=32'h00000000;
        mem[176]<=32'h00000000;
        mem[177]<=32'h00000000;
        mem[178]<=32'h00000000;
        mem[179]<=32'h00000000;
        mem[180]<=32'h00000000;
        mem[181]<=32'h00000000;
        mem[182]<=32'h00000000;
        mem[183]<=32'h00000000;
        mem[184]<=32'h00000000;
        mem[185]<=32'h00000000;
        mem[186]<=32'h00000000;
        mem[187]<=32'h00000000;
        mem[188]<=32'h00000000;
        mem[189]<=32'h00000000;
        mem[190]<=32'h00000000;
        mem[191]<=32'h00000000;
        mem[192]<=32'h00000000;
        mem[193]<=32'h00000000;
        mem[194]<=32'h00000000;
        mem[195]<=32'h00000000;
        mem[196]<=32'h00000000;
        mem[197]<=32'h00000000;
        mem[198]<=32'h00000000;
        mem[199]<=32'h00000000;
        mem[200]<=32'h00000000;
        mem[201]<=32'h00000000;
        mem[202]<=32'h00000000;
        mem[203]<=32'h00000000;
        mem[204]<=32'h00000000;
        mem[205]<=32'h00000000;
        mem[206]<=32'h00000000;
        mem[207]<=32'h00000000;
        mem[208]<=32'h00000000;
        mem[209]<=32'h00000000;
        mem[210]<=32'h00000000;
        mem[211]<=32'h00000000;
        mem[212]<=32'h00000000;
        mem[213]<=32'h00000000;
        mem[214]<=32'h00000000;
        mem[215]<=32'h00000000;
        mem[216]<=32'h00000000;
        mem[217]<=32'h00000000;
        mem[218]<=32'h00000000;
        mem[219]<=32'h00000000;
        mem[220]<=32'h00000000;
        mem[221]<=32'h00000000;
        mem[222]<=32'h00000000;
        mem[223]<=32'h00000000;
        mem[224]<=32'h00000000;
        mem[225]<=32'h00000000;
        mem[226]<=32'h00000000;
        mem[227]<=32'h00000000;
        mem[228]<=32'h00000000;
        mem[229]<=32'h00000000;
        mem[230]<=32'h00000000;
        mem[231]<=32'h00000000;
        mem[232]<=32'h00000000;
        mem[233]<=32'h00000000;
        mem[234]<=32'h00000000;
        mem[235]<=32'h00000000;
        mem[236]<=32'h00000000;
        mem[237]<=32'h00000000;
        mem[238]<=32'h00000000;
        mem[239]<=32'h00000000;
        mem[240]<=32'h00000000;
        mem[241]<=32'h00000000;
        mem[242]<=32'h00000000;
        mem[243]<=32'h00000000;
        mem[244]<=32'h00000000;
        mem[245]<=32'h00000000;
        mem[246]<=32'h00000000;
        mem[247]<=32'h00000000;
        mem[248]<=32'h00000000;
        mem[249]<=32'h00000000;
        mem[250]<=32'h00000000;
        mem[251]<=32'h00000000;
        mem[252]<=32'h00000000;
        mem[253]<=32'h00000000;
        mem[254]<=32'h00000000;
        mem[255]<=32'h00000000;
    end
    initial begin
        #10;
        $readmemh("D:/PipelineCPU/test/imem.txt",mem);
    end
    
endmodule