module WriteMem();


endmodule