module Execute();


endmodule