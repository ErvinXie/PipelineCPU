module Forwarding(
    input 

  
);




endmodule