module CPU(
    input clk,
    input rst
);
    wire[31:0] new_pc,pc;


    FetchInst(
        clk,
        rst,
        

    );






endmodule